module gate(A,Y);

    input A;
    output Y;


    not (Y,A);

endmodule